library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity {{cookiecutter.project_name}} is
  
end {{cookiecutter.project_name}};

architecture rtl of {{cookiecutter.project_name}} is
  
begin
  
end rtl;
